module and_gate(a,b,y);
	input a,b;
	output y;

	wire a,b,y;

	assign y=a&b;
endmodule
